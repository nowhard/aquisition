library verilog;
use verilog.vl_types.all;
entity logic_tb is
end logic_tb;

library verilog;
use verilog.vl_types.all;
entity sin_gen_tb is
end sin_gen_tb;
